library verilog;
use verilog.vl_types.all;
entity LFSR_vlg_vec_tst is
end LFSR_vlg_vec_tst;
