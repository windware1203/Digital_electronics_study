library verilog;
use verilog.vl_types.all;
entity p0606 is
    port(
        inputer         : in     vl_logic_vector(0 to 3);
        outputer        : out    vl_logic_vector(0 to 6)
    );
end p0606;
