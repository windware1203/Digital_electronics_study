library verilog;
use verilog.vl_types.all;
entity final is
    port(
        o1              : out    vl_logic;
        pin_name1       : in     vl_logic;
        pin_name2       : in     vl_logic;
        pin_name3       : in     vl_logic;
        pin_name4       : in     vl_logic;
        pin_name5       : in     vl_logic;
        pin_name6       : in     vl_logic;
        o2              : out    vl_logic;
        o3              : out    vl_logic;
        o4              : out    vl_logic;
        o5              : out    vl_logic;
        o6              : out    vl_logic
    );
end final;
