library verilog;
use verilog.vl_types.all;
entity final_vlg_check_tst is
    port(
        o1              : in     vl_logic;
        o2              : in     vl_logic;
        o3              : in     vl_logic;
        o4              : in     vl_logic;
        o5              : in     vl_logic;
        o6              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end final_vlg_check_tst;
