library verilog;
use verilog.vl_types.all;
entity p0606_vlg_vec_tst is
end p0606_vlg_vec_tst;
