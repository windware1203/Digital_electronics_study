library verilog;
use verilog.vl_types.all;
entity lfsr_vlg_vec_tst is
end lfsr_vlg_vec_tst;
