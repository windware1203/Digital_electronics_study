library verilog;
use verilog.vl_types.all;
entity cardNum_vlg_vec_tst is
end cardNum_vlg_vec_tst;
