library verilog;
use verilog.vl_types.all;
entity SevenStop_vlg_vec_tst is
end SevenStop_vlg_vec_tst;
